--------------------------------------------------------------------------------
-- mcu80_pkg.vhdl -- Support package for Light8080 MCU.
--
-- Contains functions used to initialize internal BRAM with object code.
--
-- This package will be used from the object code package where the program
-- initialized RAM constant is defined. If you use script obj2hdl it will 
-- take care of this for you.
-- The package is used in entity mcu80 too, and nowhere else.
--
-- Please see the LICENSE file in the project root for license matters.
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package mcu80_pkg is

-- Global signals for the TB to use in lieu of hierarchical names.
signal mon_addr :       std_logic_vector(15 downto 0);
signal mon_fetch :      std_logic;

-- Basic array type for the declaration of initialization constants.
-- This type is meant to be used to declare a constant with the object code
-- that is to be preprogrammed in an initialized RAM.
type obj_code_t is array(integer range <>) of std_logic_vector(7 downto 0);

-- Basic array type for the definition of initialized RAMs.
type ram_t is array(integer range <>) of std_logic_vector(7 downto 0);

-- Builds BRAM initialization constant from a constant CONSTRAINED byte array
-- containing the application object code.
-- The object code is placed at the beginning of the BRAM and the rest is
-- filled with zeros.
-- CAN BE USED IN SYNTHESIZABLE CODE to compute a BRAM initialization constant 
-- from a constant argument.
-- 
-- oC: Object code table (as generated by utility script obj2hdl for instance).
-- size: Size of the target memory.
-- Returns ram_t value size-bytes long, suitable for synth-time initialization 
-- of a BRAM.
function objcode_to_bram(oC : obj_code_t; size : integer) return ram_t;

-- Compute log2(A), rounding up. 
-- Use this to get the minimum width of the address bus necessary to
-- address A locations.
function log2(A : natural) return natural;

end package;

package body mcu80_pkg is

-- Builds BRAM initialization constant from a constant CONSTRAINED byte array
-- containing the application object code.
function objcode_to_bram(oC : obj_code_t; size : integer) return ram_t is
variable br : ram_t(integer range 0 to size-1);
variable i : integer;
variable obj_size : integer;
begin
    
    -- If the object code table is longer than the array size, truncate code
    if oC'length > size then
        obj_size := size;
    else
        obj_size := oC'length;
    end if;

    -- Copy object code to start of BRAM...
    for i in 0 to obj_size-1 loop
        br(i) := oC(oC'low + i);
    end loop;
    
    -- ... and fill the rest with zeros
    br(obj_size to size-1) := (others => x"00");
    
    return br;
end function objcode_to_bram;


function log2(A : natural) return natural is
begin
    for I in 1 to 30 loop -- Works for up to 32 bit integers
        if(2**I >= A) then 
            return(I);
        end if;
    end loop;
    return(30);
end function log2;

end package body;
